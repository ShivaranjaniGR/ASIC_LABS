`timescale 1 ns / 1nsmodule fa_asic1_tb3;reg a,b,c,clk;wire s,cout;fa_asic1 uut1(cout,s,a,b,c,clk);initial clk=0;initialbegin a=0;b=0;c=0;#10 a=0;b=0;c=1;#10 a=0;b=1;c=0;#10 a=0;b=1;c=1;#200 $finish;endinitialbegin$dumpfile ("fa_asic1_tb3.vcd");$dumpvars (0, fa_asic1_tb3);endalways #5 clk =~clk;endmodule